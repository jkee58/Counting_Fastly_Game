library verilog;
use verilog.vl_types.all;
entity Click_Game_tb is
end Click_Game_tb;
